library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;        -- for addition & counting
use ieee.numeric_std.all;               -- for type conversions

package Common is
	type BitMatrix is array(natural range<>,natural range<>) of std_ulogic_vector;
end Common;

package body Common is
end Common;
